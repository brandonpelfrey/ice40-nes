// Implementation of the RP2A03, which is a CPU by Ricoh combining
// the MOS 6502 (without decimal mode) and audio generation.

module mod_2a03(
  input in_2a03_clk // Clocks the CPU and APU
);

// This module mostly serves to separate APU complexity from CPU complexity.

// TODO : Wire in APU
// TODO : Wire in CPU

endmodule
