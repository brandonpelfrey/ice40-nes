// An implementation of the MOS 6502

module mod_6502(
  input in_clk_cpu
);

/// TODO : Doesn't do much yet!

endmodule
